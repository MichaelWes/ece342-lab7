package definesPkg;
   // TODO: Determine the right width
   parameter IF_ID_WIDTH = 32;
   
   // TODO: Determine the right width
   parameter ID_EX_WIDTH = 96;
   
   //TODO: Determine the right width
   parameter EX_WB_WIDTH = 96;
endpackage
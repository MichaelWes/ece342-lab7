module datapath_RF_Read
(
	clk,
	reset
);

	input clk;
	input reset;

endmodule
import definesPkg::*;

module datapath_execute
(
   clk,
   reset,
   ID_EX,
   EX_WB,
	ALUop,
	ALUop1,
	ALUop2,
	ALUout,
   o_ldst_addr,
   o_ldst_rd,
   o_ldst_wr,
   o_ldst_wrdata,
	dataw,
	regw
);
   input clk;
   input reset;   
   
   input [ID_EX_WIDTH-1:0] ID_EX;
   output logic [EX_WB_WIDTH-1:0] EX_WB;
		
	// Reassign names to ID_EX sub ranges within this module
   wire [15:0] PC;
   wire [15:0] instr;
   wire [15:0] data1; //[Rx]
   wire [15:0] data2; //[Ry]
   wire [15:0] s_ext_imm8;
   wire [15:0] s_ext_imm11;
   wire valid;
	wire [2:0] Rx;
	wire [2:0] Ry;
	wire Rx_valid, Ry_valid;
	
   assign {Rx_valid, Ry_valid, Rx, Ry, valid, s_ext_imm8, s_ext_imm11, data1, data2, PC, instr} = ID_EX;
   	
   // ALU
   output logic [2:0] ALUop;	
   output logic [15:0] ALUop1;
   output logic [15:0] ALUop2;
	input [15:0] ALUout;
	
	// ld/st signals 
	output logic [15:0] o_ldst_addr;
   output logic o_ldst_rd;
   output logic o_ldst_wr;
   output logic [15:0] o_ldst_wrdata;
	
	wire [4:0] opcode = instr[4:0];
	
	// forwarded signals from WB stage
	input [15:0] dataw;
	input [2:0] regw;
	
	// forwarded operands, or operands read from ID_EX, whichever is more recent
	logic [15:0] operand1;
	logic [15:0] operand2;
	
		// Operand forwarding logic
	always_comb begin
		operand1 = data1;
		operand2 = data2;
		if((regw == Rx) & Rx_valid) begin
			operand1 = dataw;
		end
		if((regw == Ry) & Ry_valid) begin
			operand2 = dataw;
		end
	end
	
	always_comb begin
		casex(opcode)
			// mv
			5'b00000: begin
				ALUop1 = '0;
				ALUop2 = operand2;
			end
			// add
			5'b00001: begin
				ALUop1 = operand1;
				ALUop2 = operand2;
			end
			// sub, cmp
			5'b0001x: begin
				ALUop1 = operand1;
				ALUop2 = operand2;
			end
			// mvi
			5'b10000: begin
				ALUop1 = '0;
				ALUop2 = s_ext_imm8;
			end
			// addi
			5'b10001: begin
				ALUop1 = operand1;
				ALUop2 = s_ext_imm8;
			end
			// subi, cmpi
			5'b1001x: begin
				ALUop1 = operand1;
				ALUop2 = s_ext_imm8;
			end
			5'b10110: begin
				ALUop1 = operand1;
				ALUop2 = instr[15:8]; // imm8
			end
			// TODO: ALU operands MUX for the rest of the instructions
			default: begin
				ALUop1 = 'x;
				ALUop2 = 'x;
			end
		endcase
	end

   always_comb begin
      // ALUop signal generated based on the instruction
      casex(opcode) 
         // mv, add, mvi, addi
         5'bx000x: ALUop = 3'b000; 
         // sub, cmp, subi, cmpi
         5'bx001x: ALUop = 3'b001;
			// mvhi
			5'b10110: ALUop = 3'b100;
			// TODO: operations for other instructions
         default: ALUop = '0;
      endcase
   end
	
	// Generate signals for loads and stores
	always_comb begin
		if(valid) begin
			case(opcode)
				// ld
				5'b00100: begin
					o_ldst_addr = operand2;
					o_ldst_rd = 1'b1;
					o_ldst_wr = 1'b0;
					o_ldst_wrdata = 'x;
				end
				// st
				5'b00101: begin
					o_ldst_addr = operand2;
					o_ldst_rd = 1'b0;
					o_ldst_wr = 1'b1;
					o_ldst_wrdata = operand1;
				end
				default: begin
					o_ldst_addr = 'x;
					o_ldst_wrdata = 'x;
					o_ldst_wr = '0;
					o_ldst_rd = '0;
				end
			endcase
		end else begin
			o_ldst_addr = 'x;
			o_ldst_wrdata = 'x;
			o_ldst_wr = '0;
			o_ldst_rd = '0;
		end
	end
   
	always_ff @(posedge clk) begin
		if(reset) begin
			EX_WB <= '0;
		end else begin
			// TODO: writing BT to EX/WB 
			// TODO: other values as needed
			if(valid)
				EX_WB <= {valid, data1, data2, ALUout, instr};
		end
	end
	
endmodule
package definesPkg;
	parameter IF_ID_WIDTH = 32;
	
	// TODO: Determine the right width
	parameter ID_EX_WIDTH = 64;
endpackage
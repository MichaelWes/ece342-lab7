package definesPkg;
   // TODO: Determine the right width
   parameter IF_ID_WIDTH = 33;
   
   // TODO: Determine the right width
   parameter ID_EX_WIDTH = 97;
   
   //TODO: Determine the right width
   parameter EX_WB_WIDTH = 97;
endpackage
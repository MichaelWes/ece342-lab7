package definesPkg;
   // TODO: Determine the right width
   parameter IF_ID_WIDTH = 32 + 1;
   
   // TODO: Determine the right width
   parameter ID_EX_WIDTH = 96 + 1 + 8;
   
   //TODO: Determine the right width
   parameter EX_WB_WIDTH = (16 * 5) + 1;
endpackage